LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY gtr16_tb IS
END ENTITY;

ARCHITECTURE testbench OF gtr16_tb IS
  COMPONENT gtr16
    PORT (
      in0, in1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
      cout : OUT STD_LOGIC
    );
  END COMPONENT;

  SIGNAL in0, in1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  SIGNAL cout : STD_LOGIC;

BEGIN
  GTR160 : gtr16 PORT MAP(in0, in1, cout);

  PROCESS
  BEGIN
    in0 <= "0011011100110011";
    in1 <= "0101010101000001";
    WAIT FOR 5 ns;
    in0 <= "1111111111111111";
    in1 <= "1111111111111110";
    WAIT FOR 5 ns;
    in0 <= "0101010101000001";
    in1 <= "0011011100110011";
    WAIT FOR 5 ns;
    in0 <= "1111111111111110";
    in1 <= "1111111111111111";
    WAIT FOR 5 ns;
    in0 <= "0000000000000000";
    in1 <= "0000000000000000";
    WAIT FOR 5 ns;
  END PROCESS;
END;