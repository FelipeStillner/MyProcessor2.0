LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY rom IS
    PORT (
        clk : IN STD_LOGIC;
        endereco : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
        dado : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE a_rom OF rom IS
    TYPE mem IS ARRAY (-64 TO 127) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
    CONSTANT conteudo_rom : mem := (
        -- caso endereco => conteudo
        0 => "0111111101000100",
        1 => "0000000100100100",
        2 => "0000000000111000",
        3 => "0000000000110000",
        4 => "0000000000111000",
        5 => "0000000100001111",
        6 => "0000000000111100",
        7 => "0000000000111000",
        8 => "0000000001010001",
        9 => "1111100100010110",
        10 => "0000001011100100",
        11 => "0000000000000000",
        12 => "0000000011111000",
        13 => "0000000001111100",
        14 => "0000000011111000",
        15 => "0000000011011100",
        16 => "0000000011011000",
        17 => "0000000011101101",
        18 => "0000000011011100",
        19 => "0000000011011000",
        20 => "0000000000010000",
        21 => "0000000001011000",
        22 => "0000000011010001",
        23 => "1111100100010110",
        24 => "0000000000000000",
        25 => "0000000011111000",
        26 => "0000000100001111",
        27 => "0000000011111100",
        28 => "0000000011111000",
        29 => "0000000000000000",
        30 => "0000000011111000",
        31 => "0000000010110100",
        32 => "0000000000011000",
        33 => "0000000010110001",
        34 => "0000001000010110",
        35 => "0001011100001110",
        36 => "0000000000000000",
        37 => "0001000100101100",
        38 => "0000000000111000",
        39 => "0111011000001111",
        40 => "0000000000111100",
        41 => "0000000000111000",
        42 => "0000000001110001",
        43 => "0000000000111100",
        44 => "0000000000011000",
        45 => "0000000000110001",
        46 => "1111101100010110",
        47 => "0000000000111000",
        48 => "0000000000001111",
        49 => "0000001100010110",
        50 => "0000000001111000",
        51 => "0000000010011100",
        52 => "0000101100001110",
        53 => "0000000000000000",
        54 => "0000000000000000",
        55 => "0000000000000000",
        
        -- abaixo: casos omissos => (zero em todos os bits)
        OTHERS => (OTHERS => '0')
    );
BEGIN
    PROCESS (clk)
    BEGIN
        IF (rising_edge(clk)) THEN
            dado <= conteudo_rom(to_integer(signed(endereco)));
        END IF;
    END PROCESS;
END ARCHITECTURE;