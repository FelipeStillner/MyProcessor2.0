LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY and16_tb IS
END ENTITY;

ARCHITECTURE testbench OF and16_tb IS
  COMPONENT and16
    PORT (
      in0, in1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
      out0 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
  END COMPONENT;

  SIGNAL in0, in1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  SIGNAL out0 : STD_LOGIC_VECTOR(15 DOWNTO 0);

BEGIN
  AND160 : and16 PORT MAP(in0, in1, out0);

  PROCESS
  BEGIN
    in0 <= "0011001100110011";
    in1 <= "0101010101010101";
    WAIT FOR 5 ns;
  END PROCESS;
END;