LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY leftshift16_tb IS
END ENTITY;

ARCHITECTURE testbench OF leftshift16_tb IS
  COMPONENT leftshift16
    PORT (
      in0, in1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
      out0 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
  END COMPONENT;

  SIGNAL in0, in1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  SIGNAL out0 : STD_LOGIC_VECTOR(15 DOWNTO 0);

BEGIN
  LFT160 : leftshift16 PORT MAP(in0, in1, out0);

  PROCESS
  BEGIN
    in0 <= "0011011100110011";
    in1 <= "0000000000000000";
    WAIT FOR 5 ns;
    in0 <= "1111111111111111";
    in1 <= "0000000000000001";
    WAIT FOR 5 ns;
    in0 <= "1111111011011100";
    in1 <= "0000000000000101";
    WAIT FOR 5 ns;
    in0 <= "0000100011001110";
    in1 <= "0000000000001111";
    WAIT FOR 5 ns;
  END PROCESS;
END;