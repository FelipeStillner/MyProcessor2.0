LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY leftshift16 IS
    PORT (
        in0, in1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        out0 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE behaviour OF leftshift16 IS
BEGIN
    out0 <= (in0) WHEN (in1 = "0000000000000000") ELSE
        (in0(14 DOWNTO 0) & "0") WHEN (in1 = "0000000000000001") ELSE
        (in0(13 DOWNTO 0) & "00") WHEN (in1 = "0000000000000010") ELSE
        (in0(12 DOWNTO 0) & "000") WHEN (in1 = "0000000000000011") ELSE
        (in0(11 DOWNTO 0) & "0000") WHEN (in1 = "0000000000000100") ELSE
        (in0(10 DOWNTO 0) & "00000") WHEN (in1 = "0000000000000101") ELSE
        (in0(9 DOWNTO 0) & "000000") WHEN (in1 = "0000000000000110") ELSE
        (in0(8 DOWNTO 0) & "0000000") WHEN (in1 = "0000000000000111") ELSE
        (in0(7 DOWNTO 0) & "00000000") WHEN (in1 = "0000000000001000") ELSE
        (in0(6 DOWNTO 0) & "000000000") WHEN (in1 = "0000000000001001") ELSE
        (in0(5 DOWNTO 0) & "0000000000") WHEN (in1 = "0000000000001010") ELSE
        (in0(4 DOWNTO 0) & "00000000000") WHEN (in1 = "0000000000001011") ELSE
        (in0(3 DOWNTO 0) & "000000000000") WHEN (in1 = "0000000000001100") ELSE
        (in0(2 DOWNTO 0) & "0000000000000") WHEN (in1 = "0000000000001101") ELSE
        (in0(1 DOWNTO 0) & "00000000000000") WHEN (in1 = "0000000000001110") ELSE
        (in0(0 DOWNTO 0) & "000000000000000") WHEN (in1 = "0000000000001111") ELSE
        "0000000000000000";
END ARCHITECTURE;